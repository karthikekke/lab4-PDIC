/u/ekke/PDIC/lab4-karthikekke/apr/work/saed32nm_rvt_1p9m.lef