/u/ekke/PDIC/lab4-karthikekke/apr/work/saed32sram.lef