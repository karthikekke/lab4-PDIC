/u/ekke/PDIC/lab4-karthikekke/cadence_cap_tech/tech.lef